/*
 *  TOPPERS/FMP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Multi-Processor
 * 
 *  Copyright (C) 2015,2016 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015-2018 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *  Copyright (C) 2019 by TOPPERS Project
 * 
 *  上記著作権者は，以下の(1)〜(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id: kernel.cdl 285 2018-03-21 02:55:49Z ertl-hiro $
 */

/*
 *		TOPPERS/FMPカーネルオブジェクト コンポーネント記述ファイル
 */

/*
 *  カーネルオブジェクトのコンポーネント化のためのヘッダファイル
 */
import_C("tecs_kernel.h");

/*
 *  タスク操作のシグニチャ（タスクコンテキスト用）
 */
signature sTaskRs {
	PLType("Result<(), itron::error::Error<itron::task::ActivateError>>")				activate(void);
	PLType("Result<(), itron::error::Error<itron::task::ActivateOnError>>")			migrateAndActivate([in] PLType("itron::processor::Processor") prcid);           // FMP3
	PLType("Result<usize, itron::error::Error<itron::task::CancelActivateAllError>>") cancelActivate(void);
	PLType("Result<(), itron::error::Error<itron::task::MigrateError>>")              migrate([in] PLType("itron::processor::Processor") prcid);                      // FMP3
	PLType("Result<itron::task::State, itron::error::Error<itron::task::StateError>>")             getTaskState(void);
	PLType("Result<(), itron::error::Error<itron::task::SetPriorityError>>")          	changePriority([in] PLType("itron::task::Priority") priority);
	PLType("itron::abi::ER")                                                                    changeSubPriority([in] uint_t subPriority);  // FMP3
	PLType("Result<itron::task::Priority, itron::error::Error<itron::task::PriorityError>>")       getPriority(void);
	PLType("Result<itron::task::Info, itron::error::Error<itron::task::InfoError>>")               refer(void);

	PLType("Result<(), itron::error::Error<itron::task::WakeError>>")                 wakeup(void);
	PLType("Result<usize, itron::error::Error<itron::task::CancelWakeAllError>>")     cancelWakeup(void);
	PLType("Result<(), itron::error::Error<itron::task::ReleaseWaitError>>")          releaseWait(void);
	PLType("Result<(), itron::error::Error<itron::task::SuspendError>>")              suspend(void);
	PLType("Result<(), itron::error::Error<itron::task::ResumeError>>")               resume(void);

	PLType("Result<(), itron::error::Error<itron::task::RaiseTerminationError>>")     raiseTerminate(void);
	PLType("Result<(), itron::error::Error<itron::task::TerminateError>>")            terminate(void);
};

/*
 *  タスクのセルタイプ
 *
 *  タスクはいずれかの保護ドメインに所属させなければならない．
 */
//[active, generate(FMPObjectPlugin, "TASK"), idx_is_id]
[active, generate(FMPObjectPlugin, "TASK")]
celltype tTaskRs {
	[inline] entry	sTaskRs	eTask;
	[inline] entry	siTask	eiTask;
	call	sTaskBody	cTaskBody;

	[inline] entry	siNotificationHandler	eiActivateNotificationHandler;
	[inline] entry	siNotificationHandler	eiWakeUpNotificationHandler;

	attr {
		[omit] ID				id = PL_EXP("TSKID_$id$");
		PLType("itron::task::TaskRef<'static>")			task_ref = PL_EXP("unsafe{itron::task::TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_$id$).unwrap())}");
		[omit] ATR		attribute = PL_EXP("TA_NULL");
		[omit] PRI		priority;
		[omit] size_t	stackSize;
		[omit] size_t	systemStackSize = 0;
						/* 0を，未定義を示す値として使っている */
	};

	/*
	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
	*/
};

/*
 *  セマフォ操作のシグニチャ（タスクコンテキスト用）
 */
signature sSemaphoreRs {
	PLType("Result<(), itron::error::Error<itron::semaphore::SignalError>>")			signal(void);
	PLType("Result<(), itron::error::Error<itron::semaphore::WaitError>>")				wait(void);
	PLType("Result<(), itron::error::Error<itron::semaphore::PollError>>")				waitPolling(void);
	PLType("Result<(), itron::error::Error<itron::semaphore::WaitTimeoutError>>")		waitTimeout([in] PLType("itron::time::Timeout") timeout);
	PLType("Result<(), itron::error::Error<itron::semaphore::InitializeError>>")		initialize(void);
	PLType("Result<itron::semaphore::Info, itron::error::Error<itron::semaphore::InfoError>>")				refer(void);
};

/*
 *  セマフォのセルタイプ
 */
[generate(FMPObjectPlugin, "SEMAPHORE")]
celltype tSemaphoreRs {
	[inline] entry	sSemaphoreRs	eSemaphore;
	[inline] entry	siSemaphore	eiSemaphore;

	[inline] entry	siNotificationHandler	eiNotificationHandler;

	attr {
		[omit]ID				id = PL_EXP("SEMID_$id$");
		PLType("itron::semaphore::SemaphoreRef<'static>")	semaphore_ref = PL_EXP("unsafe{itron::semaphore::SemaphoreRef::from_raw_nonnull(NonZeroI32::new(SEMID_$id$).unwrap())}");
		[omit] ATR		attribute = PL_EXP("TA_NULL");
		[omit] uint_t	initialCount;
		[omit] uint_t	maxCount = 1;
	};

	/*
	FACTORY {
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
	*/
};

/*
 *  データキュー操作のシグニチャ（タスクコンテキスト用）
 */
signature sDataqueueRs {
	PLType("Result<(), itron::error::Error<itron::dataqueue::SendError>>") 						send([in] PLType("itron::dataqueue::DataElement") data);
	PLType("Result<(), itron::error::Error<itron::dataqueue::TrySendError>>") 					sendPolling([in] PLType("itron::dataqueue::DataElement") data);
	PLType("Result<(), itron::error::Error<itron::dataqueue::SendTimeoutError>>") 				sendTimeout([in] PLType("itron::dataqueue::DataElement") data, [in] PLType("itron::time::Timeout") timeout);
	PLType("Result<(), itron::error::Error<itron::dataqueue::SendForcedError>>") 				sendForce([in] PLType("itron::dataqueue::DataElement") data);
	PLType("Result<itron::dataqueue::DataElement, itron::error::Error<itron::dataqueue::RecvError>>") 				receive(void);
	PLType("Result<itron::dataqueue::DataElement, itron::error::Error<itron::dataqueue::TryRecvError>>") 			receivePolling(void);
	PLType("Result<itron::dataqueue::DataElement, itron::error::Error<itron::dataqueue::RecvTimeoutError>>") 		receiveTimeout([in] PLType("itron::time::Timeout") timeout);
	PLType("Result<(), itron::error::Error<itron::dataqueue::InitializeError>>") 				initialize(void);
	PLType("Result<itron::dataqueue::Info, itron::error::Error<itron::dataqueue::InfoError>>")						refer(void);
};

/*
 *  データキュー操作のシグニチャ（非タスクコンテキスト用）
 */
[context("non-task")]
signature siDataqueueRs {
	PLType("Result<(), itron::error::Error<itron::dataqueue::TrySendError>>") 			sendPolling([in] PLType("itron::dataqueue::DataElement") data);
	PLType("Result<(), itron::error::Error<itron::dataqueue::SendForcedError>>") 		sendForce([in] PLType("itron::dataqueue::DataElement") data);
};

/*
 *  データキューのセルタイプ
 */
[generate(FMPObjectPlugin, "DATAQUEUE")]
celltype tDataqueueRs {
	[inline] entry	sDataqueueRs	eDataqueue;
	[inline] entry	siDataqueueRs	eiDataqueue;

	[inline] entry	siNotificationHandler	eiNotificationHandler;

	attr {
		[omit] ID				id = PL_EXP("DTQID_$id$");
		PLType("itron::dataqueue::DataqueueRef<'static>")	dataqueue_ref = PL_EXP("unsafe{itron::dataqueue::DataqueueRef::from_raw_nonnull(NonZeroI32::new(SEMID_$id$).unwrap())}");
		[omit] ATR		attribute = PL_EXP("TA_NULL");
		[omit] uint_t	dataCount = 1;
		[omit] void		*dataqueueManagementBuffer = PL_EXP("NULL");
	};

	/*
	FACTORY {
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
	*/
};


// TODO: 割込みは itron_rs で実装されていないため、暫定的な実装を行う
/*
 *  割込み要求ライン操作のシグニチャ（タスクコンテキスト用）
 */
signature sInterruptRequestRs {
	PLType("Result<(), itron::abi::ER>")		disable(void);
	PLType("Result<(), itron::abi::ER>")		enable(void);
	PLType("Result<(), itron::abi::ER>")		clear(void);
	PLType("Result<(), itron::abi::ER>")		raise(void);
	PLType("Result<bool, itron::abi::ER>")		probe(void);
};

/*
 *  割込み要求ラインのセルタイプ
 *
 *  割込み要求ラインはカーネルドメインに所属させなければならない．
 */
[active, generate(FMPHandlerPlugin, "INT_REQUEST")]
celltype tInterruptRequestRs {
	[inline] entry	sInterruptRequestRs	eInterruptRequest;

	attr {
		INTNO			interruptNumber;
		[omit] ATR		attribute = PL_EXP("TA_NULL");
		[omit] PRI		interruptPriority;
	};

	/* 警告メッセージを抑止するための記述 */
	/*
	factory {
		write("tecsgen.cfg", "");
	};
	*/
};

/*
 *  割込みサービスルーチンのセルタイプ
 *
 */
[active, generate(FMPHandlerPlugin, "INT_SERVICE_ROUTINE")]
celltype tIsrRs {
	call	siHandlerBody	ciIsrBody;

	attr {
		ID				id = PL_EXP("ISRID_$id$");
		[omit] ATR		attribute = PL_EXP("TA_NULL");
		[omit] INTNO	interruptNumber;
		[omit] PRI		isrPriority = 1;
	};

	/*
	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
		write("$ct$_factory.h", "#include \"kernel_cfg.h\"");
	};
	*/
};


/*
 *  初期化ルーチンのセルタイプ
 *
 *  初期化ルーチンはカーネルドメインに所属させなければならない．
 */
[active, generate(FMPHandlerPlugin, "INIT_ROUTINE")]
celltype tInitializeRoutineRs {
	call	sRoutineBody	cInitializeRoutineBody;

	attr {
		[omit] ATR		attribute = PL_EXP("TA_NULL");
	};

	/*
	FACTORY {
		write("tecsgen.cfg", "#include \"$ct$_tecsgen.h\"");
	};
	*/
};