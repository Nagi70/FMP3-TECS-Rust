/*
 *  カーネルオブジェクトの定義
 */
import(<kernel.cdl>);
import(<kernel_rs.cdl>);
//import("target.cdl");
import( <target_class.cdl> );

/*
 *  ターゲット非依存のセルタイプの定義
 */
import("syssvc/tSerialPort.cdl");
import("syssvc/tSerialAdapter.cdl");
import("syssvc/tSysLog.cdl");
import("syssvc/tSysLogAdapter.cdl");
import("syssvc/tLogTask.cdl");
import("syssvc/tBanner.cdl");

/*
 *  ターゲット依存部の取り込み
 */
import("target.cdl");

region rProcessor1Migratable {
   /*
    *		システムログ機能のアダプタの組上げ記述
    *
    *  システムログ機能のアダプタは，C言語で記述されたコードから，TECSベー
    *  スのシステムログ機能を呼び出すためのセルである．システムログ機能の
    *  サービスコール（syslog，syslog_0〜syslog_5，t_perrorを含む）を呼び
    *  出さない場合には，以下のセルの組上げ記述を削除してよい．
    */
   cell tSysLogAdapter SysLogAdapter {
     cSysLog = SysLog.eSysLog;
   };

   /*
    *		シリアルインタフェースドライバのアダプタの組上げ記述
    *
    *  シリアルインタフェースドライバのアダプタは，C言語で記述されたコー
    *  ドから，TECSベースのシリアルインタフェースドライバを呼び出すための
    *  セルである．シリアルインタフェースドライバのサービスコールを呼び出
    *  さない場合には，以下のセルの組上げ記述を削除してよい．
    */
   cell tSerialAdapter SerialAdapter {
     cSerialPort[0] = SerialPort1.eSerialPort;
   };

   /*
    *		システムログ機能の組上げ記述
    *
    *  システムログ機能を外す場合には，以下のセルの組上げ記述を削除し，コ
    *  ンパイルオプションに-DTOPPERS_OMIT_SYSLOGを追加すればよい．ただし，
    *  システムログタスクはシステムログ機能を使用するため，それも外すこと
    *  が必要である．また，システムログ機能のアダプタも外さなければならな
    *  い．tecsgenが警告メッセージを出すが，無視してよい．
    */
   cell tSysLog SysLog {
     logBufferSize = 32;					/* ログバッファのサイズ */
     initLogMask = C_EXP("LOG_UPTO(LOG_NOTICE)");
                       /* ログバッファに記録すべき重要度 */
     initLowMask = C_EXP("LOG_UPTO(LOG_EMERG)");
                         /* 低レベル出力すべき重要度 */
     /* 低レベル出力との結合 */
     cPutLog = PutLogTarget.ePutLog;
   };

   /*
    *		シリアルインタフェースドライバの組上げ記述
    *
    *  シリアルインタフェースドライバを外す場合には，以下のセルの組上げ記
    *  述を削除すればよい．ただし，システムログタスクはシリアルインタフェー
    *  スドライバを使用するため，それも外すことが必要である．また，シリア
    *  ルインタフェースドライバのアダプタも外さなければならない．
    */
   cell tSerialPort SerialPort1 {
     receiveBufferSize = 256;			/* 受信バッファのサイズ */
     sendBufferSize    = 256;			/* 送信バッファのサイズ */

     /* ターゲット依存部との結合 */
     cSIOPort = SIOPortTarget1.eSIOPort;
     eiSIOCBR <= SIOPortTarget1.ciSIOCBR;	/* コールバック */
   };

   /*
    *		システムログタスクの組上げ記述
    *
    *  システムログタスクを外す場合には，以下のセルの組上げ記述を削除すれ
    *  ばよい．
    */
   cell tLogTask LogTask {
     priority  = 3;					/* システムログタスクの優先度 */
     stackSize = LogTaskStackSize;	/* システムログタスクのスタックサイズ */

     /* シリアルインタフェースドライバとの結合 */
     cSerialPort        = SerialPort1.eSerialPort;
     cnSerialPortManage = SerialPort1.enSerialPortManage;

     /* システムログ機能との結合 */
     cSysLog = SysLog.eSysLog;

     /* 低レベル出力との結合 */
     cPutLog = PutLogTarget.ePutLog;
   };

   /*
    *		カーネル起動メッセージ出力の組上げ記述
    *
    *  カーネル起動メッセージの出力を外す場合には，以下のセルの組上げ記述
    *  を削除すればよい．
    */
   cell tBanner Banner {
     /* 属性の設定 */
     targetName      = BannerTargetName;
     copyrightNotice = BannerCopyrightNotice;
   };
};

celltype tMeasure {
  call sTaskRs cTask;
  call sTaskRs cTaskmig;
  call sSemaphoreRs cSemaphore;
  entry sTaskBody eTaskbody;
};

celltype tReset {
  call sTaskRs cTask;
  call sTaskRs cTaskself;
  call sTaskRs cTaskmig;
  call sSemaphoreRs cSemaphore;
  entry sTaskBody eReset;
};

celltype tTaskbodyRs2 {
  entry sTaskBody eTaskbody;
};

celltype tSelfReset {
  call sTaskRs cTaskself;
  entry sTaskBody eSelfReset;
  call sSemaphoreRs cSemaphore;
};

[class(FMP,"CLS_PRC1")]
region rProcessor1Symmetric{

    [generate(RustFMP3Plugin, "TASK, lib")]
    cell tTaskRs Task1_1 {
        /* 呼び口の結合 */
        cTaskBody = rProcessor1Symmetric::Measure.eTaskbody;
        /* 属性の設定 */
        id = C_EXP("TSKID_1_1");
        task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_1_1).unwrap())}");
        priority = 7;
        stackSize = 2048;
        attribute = C_EXP("TA_ACT");
    };

    [generate (RustFMP3Plugin, "lib")]
    cell tMeasure Measure {
      cTask = rProcessor2Symmetric::Task2_2.eTask;
      cTaskmig = rProcessorAllMig::Taskmig.eTask;
      cSemaphore = rProcessorAllMig::Semaphore.eSemaphore;
    };
};

[class(FMP,"CLS_ALL_PRC1")]
region rProcessorAllMig{
    [generate (RustFMP3Plugin, "SEMAPHORE, lib")]
    cell tSemaphoreRs Semaphore {
      id = C_EXP("SEMID_1");
      semaphore_ref = C_EXP("unsafe{SemaphoreRef::from_raw_nonnull(NonZeroI32::new(SEMID_1).unwrap())}");
      initialCount = 1;
    };

    [generate(RustFMP3Plugin, "TASK, lib")]
    cell tTaskRs Taskmig {
        /* 呼び口の結合 */
        cTaskBody = rProcessorAllMig::Taskbody1_2.eTaskbody;
        /* 属性の設定 */
        id = C_EXP("TSKID_MIG");
        task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_MIG).unwrap())}");
        priority = 10;
        stackSize = 2048;
        attribute = C_EXP("TA_ACT");
    };

    [generate (RustFMP3Plugin, "lib")]
    cell tTaskbodyRs2 Taskbody1_2 {
    };
};

[class(FMP,"CLS_PRC2")]
region rProcessor2Symmetric{

    [generate(RustFMP3Plugin, "TASK, lib")]
    cell tTaskRs Task2_1 {
        /* 呼び口の結合 */
        cTaskBody = rProcessor2Symmetric::Reset.eReset;
        /* 属性の設定 */
        id = C_EXP("TSKID_2_1");
        task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_2_1).unwrap())}");
        priority = 7;
        stackSize = 2048;
        attribute = C_EXP("TA_ACT");
    };

    [generate (RustFMP3Plugin, "lib")]
    cell tReset Reset {
      cTask = rProcessor2Symmetric::Task2_2.eTask;
      cTaskself = rProcessor2Symmetric::Task2_1.eTask;
      cTaskmig = rProcessorAllMig::Taskmig.eTask;
      cSemaphore = rProcessorAllMig::Semaphore.eSemaphore;
    };

    [generate(RustFMP3Plugin, "TASK, lib")]
    cell tTaskRs Task2_2 {
        /* 呼び口の結合 */
        cTaskBody = rProcessor2Symmetric::SelfReset.eSelfReset;
        /* 属性の設定 */
        id = C_EXP("TSKID_2_2");
        task_ref = C_EXP("unsafe{TaskRef::from_raw_nonnull(NonZeroI32::new(TSKID_2_2).unwrap())}");
        priority = 10;
        stackSize = 2048;
        attribute = C_EXP("TA_NULL");
    };

    [generate (RustFMP3Plugin, "lib")]
    cell tSelfReset SelfReset {
      cTaskself = rProcessor2Symmetric::Task2_2.eTask;
      cSemaphore = rProcessorAllMig::Semaphore.eSemaphore;
    };
};



